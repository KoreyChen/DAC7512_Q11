library verilog;
use verilog.vl_types.all;
entity dac7512_vlg_tst is
    generic(
        clk_set         : integer := 20
    );
end dac7512_vlg_tst;
